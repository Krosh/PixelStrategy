name:Country
infantry:0
size:859
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:1910
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:1961
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:1472
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:976
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:2684
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:383
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:2331
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:1464
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:2044
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:1056
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:1549
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:1631
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:1265
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:1457
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:3633
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:5893
peons:150
grow:0
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:2870
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:2925
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
name:Country
infantry:0
size:1637
peons:150
grow:0
food:200
money:100
artillery:0
scientists:100
cavalry:0
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
research
name:Research
endValue:100
curValue:60
level:1
scientistsCount:10
end
